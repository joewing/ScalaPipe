
module ap_addI(a_in, b_in, c_out);

   parameter WIDTH = 32;
   input wire [WIDTH-1:0] a_in;
   input wire [WIDTH-1:0] b_in;
   output wire [WIDTH-1:0] c_out;

   assign c_out = a_in + b_in;

endmodule

module ap_subI(a_in, b_in, c_out);

   parameter WIDTH = 32;
   input wire [WIDTH-1:0] a_in;
   input wire [WIDTH-1:0] b_in;
   output wire [WIDTH-1:0] c_out;

   assign c_out = a_in - b_in;

endmodule

